library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.common.all;

entity imem is
    port(
        addr : in std_logic_vector(5 downto 0);
        dout : out word);
end  imem;

architecture behavioral of imem is
type rom_arr is array(0 to 55) of word;

constant mem:rom_arr:=
    (
     --              	nprimes:
     --
    x"00300793", --  0 0000 93073000 		  0000 0000 0011 0000 0000 0111 1 0010011   li	    a5,3
    x"00050613", --  1 0004 13060500 		  000000000000 01010 000 01100 0010011      mv	    a2,a0
    x"08A7FC63", --  2 0008 63FCA708 		  0 000100 01010 01111 111 1100 0 1100011   bleu	  a0,a5,.L2
    x"000005B7", --  3 000c B7050000 		  0000 0000 0000 0000 0000 0101 1011 0111   lui	    a1,%hi(testarray+8)
    x"00000337", --  4 0010 37030000      0000 0000 0000 0000 0000 0011 0011 0111   lui	    t1,%hi(testarray)
    x"00858513", --  5 0014 13858500 		  0000 0000 1000 0101 1000 0101 0001 0011   addi    a0,a1,%lo(testarray+8)
    x"00200693", --  6 0018 93062000 		  0000 0000 0010 0000 0000 0110 1001 0011   li	    a3,2
    x"00858593", --  7 001c 93858500 		  0000 0000 1000 0101 1000 0101 1001 0011   addi	  a1,a1,%lo(testarray+8)
    x"00030313", --  8 0020 13030300 		  0000 0000 0000 0011 0000 0011 0001 0011   addi	  t1,t1,%lo(testarray)
    x"00100893", --  9 0024 93081000 		  0000 0000 0001 0000 0000 1000 1001 0011   li	    a7,1
    x"0140006F", -- 10 0028 6F004001 		  0000 0001 0100 0000 0000 0000 0 1101111   j	      .L5
    --                               	.L3:
    x"00168693", -- 11 002c 93861600 		  0000 0000 0001 0110 1000 0110 1001 0011   addi	  a3,a3,1
    x"02D687B3", -- 12 0030 B387D602 		  0000 0010 1101 0110 1000 0111 1011 0011   mul	    a5,a3,a3
    x"00458593", -- 13 0034 93854500 		  0000 0000 0100 0101 1000 0101 1001 0011   addi	  a1,a1,4
    x"04F66063", -- 14 0038 6360F604 		  0 0000100 1111 01100 110 0000 0 1100011   bgtu	  a5,a2,.L7
    --              	                .L5:
    x"0005A783", -- 15 003c 83A70500 		  0000 0000 0000 0101 1010 0111 1000 0011   lw	    a5,0(a1)
    x"FE0796E3", -- 16 0040 E39607FE 		  1 111111 00000 01111 001 0110 1 1100011   bnez	  a5,.L3
    x"00169713", -- 17 0044 13971600 		  0000 0000 0001 0110 1001 0111 0001 0011   slli	  a4,a3,1
    x"FEE662E3", -- 18 0048 E362E6FE 		  1 111111 01110 01100 110 0010 1 1100011   bltu	  a2,a4,.L3
    x"00369793", -- 19 004c 93973600 		  0000 0000 0011 0110 1001 0111 1001 0011   slli	  a5,a3,3
    x"00269813", -- 20 0050 13982600 		  0000 0000 0010 0110 1001 1000 0001 0011   slli	  a6,a3,2
    x"006787B3", -- 21 0054 B3876700 		  0000 0000 0110 0111 1000 0111 1011 0011   add	    a5,a5,t1
    --              	                .L4:
    x"0117A023", -- 22 0058 23A01701 		  0000 0001 0001 0111 1010 0000 0010 0011   sw	    a7,0(a5)
    x"00D70733", -- 23 005c 3307D700 		  0000 0000 1101 0111 0000 0111 0011 0011   add	    a4,a4,a3
    x"010787B3", -- 24 0060 B3870701 		  0000 0001 0000 0111 1000 0111 1011 0011   add	    a5,a5,a6
    x"FEE67AE3", -- 25 0064 E37AE6FE 		  1 111111 01110 01100 111 1010 1 1100011   bgeu	  a2,a4,.L4
    x"00168693", -- 26 0068 93861600 		  0000 0000 0001 0110 1000 0110 1001 0011   addi	  a3,a3,1
    x"02D687B3", -- 27 006c B387D602 		  0000 0010 1101 0110 1000 0111 1011 0011   mul	    a5,a3,a3
    x"00458593", -- 28 0070 93854500 		  0000 0000 0100 0101 1000 0101 1001 0011   addi	  a1,a1,4
    x"FCF674E3", -- 29 0074 E374F6FC 		  1 111110 01111 01100 111 0100 1 1100011   bleu	  a5,a2,.L5
    --                               	.L7:
    x"00050713", -- 30 0078 13070500 		  0000 0000 0000 0101 0000 0111 0001 0011   mv	    a4,a0
    x"00200693", -- 31 007c 93062000 		  0000 0000 0010 0000 0000 0110 1001 0011   li	    a3,2
    x"00000513", -- 32 0080 13050000 		  0000 0000 0000 0000 0000 0101 0001 0011   li	    a0,0
    --                              	.L6:
    x"00072783", -- 33 0084 83270700 		  0000 0000 0000 0111 0010 0111 1000 0011   lw	    a5,0(a4)
    x"00168693", -- 34 0088 93861600 		  0000 0000 0001 0110 1000 0110 1001 0011   addi	  a3,a3,1
    x"00470713", -- 35 008c 13074700 		  0000 0000 0100 0111 0000 0111 0001 0011   addi	  a4,a4,4
    x"0017B793", -- 36 0090 93B71700 		  0000 0000 0001 0111 1011 0111 1001 0011   seqz	  a5,a5
    x"00F50533", -- 37 0094 3305F500 		  0000 0000 1111 0101 0000 0101 0011 0011   add	    a0,a0,a5
    x"FED676E3", -- 38 0098 E376D6FE 		  1 111111 01101 01100 111 0110 1 1100011  	bleu    a3,a2,.L6
    x"00008067", -- 39 009c 67800000 		  0000 0000 0000 0000 1000 0000 0 1100111   ret
    --                               	.L2:
    x"00100793", -- 40 00a0 93071000 		  0000 0000 0001 0000 0000 0111 1001 0011   li	    a5,1
    x"00A7E663", -- 41 00a4 63E6A700 		  0 000000 01010 01111 110 0110 0 1100011   bgtu	  a0,a5,.L16
    x"00000513", -- 42 00a8 13050000 		  0000 0000 0000 0000 0000 0101 0001 0011   li	    a0,0
    x"00008067", -- 43 00ac 67800000 		  0000 0000 0000 0000 1000 0000 0 1100111   ret
    --
    --               	.L16:
    x"00000737", -- 45 00b0 37070000 	    0000 0000 0000 0000 0000 0111 0011 0111  lui	a4,%hi(testarray+8)
    x"00870513", -- 46 00b4 13058700 		  0000 0000 1000 0111 0000 0101 0001 0011  addi	a0,a4,%lo(testarray+8)
    x"FC1FF06F", -- 47 00b8 6FF01FFC 		  1 1111100 000 1 11111111 00000 1101111   j	.L7
    --
    --                              	main:
    --
    x"FF010113", -- 48 0000 130101FF 		1111 1111 0000 0001 0000 00010 0010011    addi	   sp,sp,-16
    x"06400513", -- 49 0004 13054006 		0000011 00100 00000 000 01010 0010011     li	     a0,100
    x"00112623", -- 50 0008 23261100 		0000000 00001 00010 010 01100 0100011     sw	     ra,12(sp)
    x"00000097", -- 51 000c 97000000 		0000 0000 0000 00000 000 00001 0010111    call	   nprimes
    x"000080E7", -- 51      E7800000    0000 0000 0000 0000  100 00000  1100111
    x"00C12083", -- 52 0014 8320C100 		0000 0000 1100 0001 0010 0000 1000 0011   lw	     ra,12(sp)
    x"00000513", -- 53 0018 13050000 		0000 0000 0000 0000 0000 0101 0001 0011   li	     a0,0
    x"01010113", -- 54 001c 13010101 		0000 0001 0000 0001 0000 0001 0001 0011   addi	   sp,sp,16
    x"00008067");-- 55 0020 67800000 		0000 0000 0000 0000 1000 00000  1100111   jr	     ra

begin
	dout<=mem(conv_integer(addr));
end behavioral;
