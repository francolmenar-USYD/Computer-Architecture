library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library work;
use work.common.all;

entity imem is
    port(
        addr : in std_logic_vector(3 downto 0);
        dout : out word);
end imem;

architecture behavioral of imem is
type rom_arr is array(0 to 15) of word;

constant mem:rom_arr:=
    (

    x"00000793", --   8 0000 93070000     1001 0011 0000 0111 0000 0000 0000 0000   li      a5,0
    x"00C00693", --   9 0004 9306C000     1001 0011 0000 0110 1100 0000 0000 0000   li      a3,12
                  --  10                    .L2:
    x"00279713", --  11 0008 13972700     0001 0011 1001 0111 0010 0111 0000 0000   sll     a4,a5,2
    x"00F72023", --  12 000c 2320F700     0010 0011 0010 0000 1111 0111 0000 0000   sw      a5,0(a4)
    x"00178793", --  13 0010 93871700     1001 0011 1000 0111 0001 0111 0000 0000   add     a5,a5,1
    x"FED79AE3", --  14 0014 E39AD7FE     1110 0011 1001 1010 1101 0111 1111 1110   bne     a5,a3,.L2
    x"00000513", --  15 0018 13050000     0001 0011 0000 0101 0000 0000 0000 0000   li      a0,0
    x"00008067", --  16 001c 67800000     0110 0111 1000 0000 0000 0000 0000 0000   ret
    x"00000013", --       13000000        0001 0011 0000 0000 0000 0000 0000 0000   nop
    x"00000013", --       13000000                nop
    x"00000013", --       13000000                nop
    x"00000013", --       13000000                nop
    x"00000013", --       13000000                nop
    x"00000013", --       13000000                nop
    x"00000013", --       13000000                nop
    x"00000013"); --      13000000                nop

     --
     -- 1              	  .file	"nprimes.c"
     -- 2              		.option nopic
     -- 3              		.text
     -- 4              		.align	2
     -- 5              		.globl	nprimes
     -- 6              		.type	nprimes, @function
     -- 7              	nprimes:
    -- x"00300793", --  8 0000 93073000 		  1001 0011 0000 0111 0011 0000 0000 0000   li	    a5,3
    -- x"00050613", --  9 0004 13060500 		  0001 0011 0000 0110 0000 0101 0000 0000   mv	    a2,a0
    -- x"08A7FC63", -- 10 0008 63FCA708 		  0110 0011 1111 1100 1010 0111 0000 1000   bleu	  a0,a5,.L2
    -- x"000005B7", -- 11 000c B7050000 		  1011 0111 0000 0101 0000 0000 0000 0000   lui	    a1,%hi(testarray+8)
    -- x"00000337", -- 12 0010 37030000      0011 0111 0000 0011 0000 0000 0000 0000   lui	    t1,%hi(testarray)
    -- x"00858513", -- 13 0014 13858500 		  0001 0011 1000 0101 1000 0101 0000 0000   addi    a0,a1,%lo(testarray+8)
    -- x"00200693", -- 14 0018 93062000 		  1001 0011 0000 0110 0010 0000 0000 0000   li	    a3,2
    -- x"00858593", -- 15 001c 93858500 		  1001 0011 1000 0101 1000 0101 0000 0000   addi	  a1,a1,%lo(testarray+8)
    -- x"00030313", -- 16 0020 13030300 		  0001 0011 0000 0011 0000 0011 0000 0000   addi	  t1,t1,%lo(testarray)
    -- x"00100893", -- 17 0024 93081000 		  1001 0011 0000 1000 0001 0000 0000 0000   li	    a7,1
    -- x"0140006F", -- 18 0028 6F004001 		  0110 1111 0000 0000 0100 0000 0000 0001   j	      .L5
    -- x"00000000", -- 19              	.L3:
    -- x"00168693", -- 20 002c 93861600 		  1001 0011 1000 0110 0001 0110 0000 0000   addi	  a3,a3,1
    -- x"02D687B3", -- 21 0030 B387D602 		  1011 0011 1000 0111 1101 0110 0000 0010   mul	    a5,a3,a3
    -- x"00458593", -- 22 0034 93854500 		  1001 0011 1000 0101 0100 0101 0000 0000   addi	  a1,a1,4
    -- x"04F66063", -- 23 0038 6360F604 		  0110 0011 0110 0000 1111 0110 0000 0100   bgtu	  a5,a2,.L7
    -- x"00000000", -- 24              	.L5:
    -- x"0005A783", -- 25 003c 83A70500 		  1000 0011 1010 0111 0000 0101 0000 0000   lw	    a5,0(a1)
    -- x"FE0796E3", -- 26 0040 E39607FE 		  1110 0011 1001 0110 0000 0111 1111 1110   bnez	  a5,.L3
    -- x"00169713", -- 27 0044 13971600 		  0001 0011 1001 0111 0001 0110 0000 0000   slli	  a4,a3,1
    -- x"FEE662E3", -- 28 0048 E362E6FE 		  1110 0011 0110 0010 1110 0110 1111 1110   bltu	  a2,a4,.L3
    -- x"00369793", -- 29 004c 93973600 		  1001 0011 1001 0111 0011 0110 0000 0000   slli	  a5,a3,3
    -- x"00269813", -- 30 0050 13982600 		  0001 0011 1001 1000 0010 0110 0000 0000   slli	  a6,a3,2
    -- x"006787B3", -- 31 0054 B3876700 		  1011 0011 1000 0111 0110 0111 0000 0000   add	    a5,a5,t1
    -- x"00000000", -- 32              	.L4:
    -- x"0117A023", -- 33 0058 23A01701 		  0010 0011 1010 0000 0001 0111 0000 0001   sw	    a7,0(a5)
    -- x"00D70733", -- 34 005c 3307D700 		  0011 0011 0000 0111 1101 0111 0000 0000   add	    a4,a4,a3
    -- x"010787B3", -- 35 0060 B3870701 		  1011 0011 1000 0111 0000 0111 0000 0001   add	    a5,a5,a6
    -- x"FEE67AE3", -- 36 0064 E37AE6FE 		  1110 0011 0111 1010 1110 0110 1111 1110   bgeu	  a2,a4,.L4
    -- x"00168693", -- 37 0068 93861600 		  1001 0011 1000 0110 0001 0110 0000 0000   addi	  a3,a3,1
    -- x"02D687B3", -- 38 006c B387D602 		  1011 0011 1000 0111 1101 0110 0000 0010   mul	    a5,a3,a3
    -- x"00458593", -- 39 0070 93854500 		  1001 0011 1000 0101 0100 0101 0000 0000   addi	  a1,a1,4
    -- x"FCF674E3", -- 40 0074 E374F6FC 		  1110 0011 0111 0100 1111 0110 1111 1100   bleu	  a5,a2,.L5
    -- x"00000000", -- 41              	.L7:
    -- x"00050713", -- 42 0078 13070500 		  0001 0011 0000 0111 0000 0101 0000 0000   mv	    a4,a0
    -- x"00200693", -- 43 007c 93062000 		  1001 0011 0000 0110 0010 0000 0000 0000   li	    a3,2
    -- x"00000513", -- 44 0080 13050000 		  0001 0011 0000 0101 0000 0000 0000 0000   li	    a0,0
    -- x"00000000", -- 45              	.L6:
    -- x"00072783", -- 46 0084 83270700 		  1000 0011 0010 0111 0000 0111 0000 0000   lw	    a5,0(a4)
    -- x"00168693", -- 47 0088 93861600 		  1001 0011 1000 0110 0001 0110 0000 0000   addi	  a3,a3,1
    -- x"00470713", -- 48 008c 13074700 		  0001 0011 0000 0111 0100 0111 0000 0000   addi	  a4,a4,4
    -- x"0017B793", -- 49 0090 93B71700 		  1001 0011 1011 0111 0001 0111 0000 0000   seqz	  a5,a5
    -- x"00F50533", -- 50 0094 3305F500 		  0011 0011 0000 0101 1111 0101 0000 0000   add	    a0,a0,a5
    -- x"FED676E3", -- 51 0098 E376D6FE 		  1110 0011 0111 0110 1101 0110 1111 1110  	bleu    a3,a2,.L6
    -- x"00008067", -- 52 009c 67800000 		  0110 0111 1000 0000 0000 0000 0000 0000   ret
    -- x"00000000", -- 53              	.L2:
    -- x"00100793", -- 54 00a0 93071000 		  1001 0011 0000 0111 0001 0000 0000 0000   li	    a5,1
    -- x"00A7E663", -- 55 00a4 63E6A700 		  0110 0011 1110 0110 1010 0111 0000 0000   bgtu	  a0,a5,.L16
    -- x"00000513", -- 56 00a8 13050000 		  0001 0011 0000 0101 0000 0000 0000 0000   li	    a0,0
    -- x"00008067", -- 57 00ac 67800000 		  0110 0111 1000 0000 0000 0000 0000 0000   ret
    --
    -- x"00000000", --     GAS LISTING nprimes.s 			page 2
    -- --
    -- --
    -- x"00000000", --   58              	.L16:
    -- x"00000737", --   59 00b0 37070000 		lui	a4,%hi(testarray+8)
    -- x"00870513", --   60 00b4 13058700 		addi	a0,a4,%lo(testarray+8)
    -- x"FC1FF06F", --   61 00b8 6FF01FFC 		j	.L7
    -- x"", --   62              		.size	nprimes, .-nprimes
    -- x"", --   63              		.section	.text.startup,'ax',@progbits
    -- x"", --   64              		.align	2
    -- x"", --   65              		.globl	main
    -- x"", --   66              		.type	main, @function
    -- x"", --   67              	main:
    -- x"FF010113", --   68 0000 130101FF 		0001 0011 0000 0001 0000 0001 1111 1111   addi	   sp,sp,-16
    -- x"06400513", --   69 0004 13054006 		0001 0011 0000 0101 0100 0000 0000 0110   li	     a0,100
    -- x"00112623", --   70 0008 23261100 		0010 0011 0010 0110 0001 0001 0000 0000   sw	     ra,12(sp)
    -- x"00000097", --   71 000c 97000000 		1001 0111 0000 0000 0000 0000 0000 0000   call	   nprimes
    -- x"000080E7", --   71      E7800000    1110 0111 1000 0000 0000 0000 0000 0000
    -- x"00C12083", --   72 0014 8320C100 		1000 0011 0010 0000 1100 0001 0000 0000   lw	     ra,12(sp)
    -- x"00000513", --   73 0018 13050000 		0001 0011 0000 0101 0000 0000 0000 0000   li	     a0,0
    -- x"01010113", --   74 001c 13010101 		0001 0011 0000 0001 0000 0001 0000 0001   addi	   sp,sp,16
    -- x"00008067", --   75 0020 67800000 		0110 0111 1000 0000 0000 0000 0000 0000   jr	     ra
    -- x"", --   76              		.size	main, .-main
    -- x"", --   77              		.comm	testarray,262140,4
    -- x"", --   78              		.ident	'GCC: (GNU) 8.1.0'
    --
    -- GAS LISTING nprimes.s 			page 3
    --
    --
    -- DEFINED SYMBOLS
    --                             *ABS*:0000000000000000 nprimes.c
    --            nprimes.s:7      .text:0000000000000000 nprimes
    --                             *COM*:000000000003fffc testarray
    --            nprimes.s:67     .text.startup:0000000000000000 main
    --            nprimes.s:53     .text:00000000000000a0 .L2
    --            nprimes.s:24     .text:000000000000003c .L5
    --            nprimes.s:41     .text:0000000000000078 .L7
    --            nprimes.s:19     .text:000000000000002c .L3
    --            nprimes.s:32     .text:0000000000000058 .L4
    --            nprimes.s:45     .text:0000000000000084 .L6
    --            nprimes.s:58     .text:00000000000000b0 .L16

begin
	dout<=mem(conv_integer(addr));
end behavioral;
